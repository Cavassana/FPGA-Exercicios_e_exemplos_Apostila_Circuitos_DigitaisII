ENTITY atividade2_item1  IS -- atrib_1
PORT ( x1	 :IN INTEGER;   -- porta entrada
		 y1, Z1:OUT INTEGER);	-- porta entrada
END;
